library ieee;
use ieee.std_logic_1164.all;
use work.aes128Pkg.all;
use IEEE.numeric_std.all;

entity mixColumn is
  
	port (
		In_DI  : in  Matrix;
		Out_DO : out Matrix);

end entity mixColumn;


-------------------------------------------------------------------------------
--! @brief Behavioral architecture of the "MixColumn" function.
-------------------------------------------------------------------------------
architecture Behavioral of mixColumn is
  
  constant times2 : ByteArray := (
	16#00#,16#02#,16#04#,16#06#,16#08#,16#0a#,16#0c#,16#0e#,16#10#,16#12#,16#14#,16#16#,16#18#,16#1a#,16#1c#,16#1e#,
	16#20#,16#22#,16#24#,16#26#,16#28#,16#2a#,16#2c#,16#2e#,16#30#,16#32#,16#34#,16#36#,16#38#,16#3a#,16#3c#,16#3e#,
	16#40#,16#42#,16#44#,16#46#,16#48#,16#4a#,16#4c#,16#4e#,16#50#,16#52#,16#54#,16#56#,16#58#,16#5a#,16#5c#,16#5e#,
	16#60#,16#62#,16#64#,16#66#,16#68#,16#6a#,16#6c#,16#6e#,16#70#,16#72#,16#74#,16#76#,16#78#,16#7a#,16#7c#,16#7e#,
	16#80#,16#82#,16#84#,16#86#,16#88#,16#8a#,16#8c#,16#8e#,16#90#,16#92#,16#94#,16#96#,16#98#,16#9a#,16#9c#,16#9e#,
	16#a0#,16#a2#,16#a4#,16#a6#,16#a8#,16#aa#,16#ac#,16#ae#,16#b0#,16#b2#,16#b4#,16#b6#,16#b8#,16#ba#,16#bc#,16#be#,
	16#c0#,16#c2#,16#c4#,16#c6#,16#c8#,16#ca#,16#cc#,16#ce#,16#d0#,16#d2#,16#d4#,16#d6#,16#d8#,16#da#,16#dc#,16#de#,
	16#e0#,16#e2#,16#e4#,16#e6#,16#e8#,16#ea#,16#ec#,16#ee#,16#f0#,16#f2#,16#f4#,16#f6#,16#f8#,16#fa#,16#fc#,16#fe#,
	16#1b#,16#19#,16#1f#,16#1d#,16#13#,16#11#,16#17#,16#15#,16#0b#,16#09#,16#0f#,16#0d#,16#03#,16#01#,16#07#,16#05#,
	16#3b#,16#39#,16#3f#,16#3d#,16#33#,16#31#,16#37#,16#35#,16#2b#,16#29#,16#2f#,16#2d#,16#23#,16#21#,16#27#,16#25#,
	16#5b#,16#59#,16#5f#,16#5d#,16#53#,16#51#,16#57#,16#55#,16#4b#,16#49#,16#4f#,16#4d#,16#43#,16#41#,16#47#,16#45#,
	16#7b#,16#79#,16#7f#,16#7d#,16#73#,16#71#,16#77#,16#75#,16#6b#,16#69#,16#6f#,16#6d#,16#63#,16#61#,16#67#,16#65#,
	16#9b#,16#99#,16#9f#,16#9d#,16#93#,16#91#,16#97#,16#95#,16#8b#,16#89#,16#8f#,16#8d#,16#83#,16#81#,16#87#,16#85#,
	16#bb#,16#b9#,16#bf#,16#bd#,16#b3#,16#b1#,16#b7#,16#b5#,16#ab#,16#a9#,16#af#,16#ad#,16#a3#,16#a1#,16#a7#,16#a5#,
	16#db#,16#d9#,16#df#,16#dd#,16#d3#,16#d1#,16#d7#,16#d5#,16#cb#,16#c9#,16#cf#,16#cd#,16#c3#,16#c1#,16#c7#,16#c5#,
	16#fb#,16#f9#,16#ff#,16#fd#,16#f3#,16#f1#,16#f7#,16#f5#,16#eb#,16#e9#,16#ef#,16#ed#,16#e3#,16#e1#,16#e7#,16#e5#);
	
constant times3 : ByteArray := (
	16#00#,16#03#,16#06#,16#05#,16#0c#,16#0f#,16#0a#,16#09#,16#18#,16#1b#,16#1e#,16#1d#,16#14#,16#17#,16#12#,16#11#,
	16#30#,16#33#,16#36#,16#35#,16#3c#,16#3f#,16#3a#,16#39#,16#28#,16#2b#,16#2e#,16#2d#,16#24#,16#27#,16#22#,16#21#,
	16#60#,16#63#,16#66#,16#65#,16#6c#,16#6f#,16#6a#,16#69#,16#78#,16#7b#,16#7e#,16#7d#,16#74#,16#77#,16#72#,16#71#,
	16#50#,16#53#,16#56#,16#55#,16#5c#,16#5f#,16#5a#,16#59#,16#48#,16#4b#,16#4e#,16#4d#,16#44#,16#47#,16#42#,16#41#,
	16#c0#,16#c3#,16#c6#,16#c5#,16#cc#,16#cf#,16#ca#,16#c9#,16#d8#,16#db#,16#de#,16#dd#,16#d4#,16#d7#,16#d2#,16#d1#,
	16#f0#,16#f3#,16#f6#,16#f5#,16#fc#,16#ff#,16#fa#,16#f9#,16#e8#,16#eb#,16#ee#,16#ed#,16#e4#,16#e7#,16#e2#,16#e1#,
	16#a0#,16#a3#,16#a6#,16#a5#,16#ac#,16#af#,16#aa#,16#a9#,16#b8#,16#bb#,16#be#,16#bd#,16#b4#,16#b7#,16#b2#,16#b1#,
	16#90#,16#93#,16#96#,16#95#,16#9c#,16#9f#,16#9a#,16#99#,16#88#,16#8b#,16#8e#,16#8d#,16#84#,16#87#,16#82#,16#81#,
	16#9b#,16#98#,16#9d#,16#9e#,16#97#,16#94#,16#91#,16#92#,16#83#,16#80#,16#85#,16#86#,16#8f#,16#8c#,16#89#,16#8a#,
	16#ab#,16#a8#,16#ad#,16#ae#,16#a7#,16#a4#,16#a1#,16#a2#,16#b3#,16#b0#,16#b5#,16#b6#,16#bf#,16#bc#,16#b9#,16#ba#,
	16#fb#,16#f8#,16#fd#,16#fe#,16#f7#,16#f4#,16#f1#,16#f2#,16#e3#,16#e0#,16#e5#,16#e6#,16#ef#,16#ec#,16#e9#,16#ea#,
	16#cb#,16#c8#,16#cd#,16#ce#,16#c7#,16#c4#,16#c1#,16#c2#,16#d3#,16#d0#,16#d5#,16#d6#,16#df#,16#dc#,16#d9#,16#da#,
	16#5b#,16#58#,16#5d#,16#5e#,16#57#,16#54#,16#51#,16#52#,16#43#,16#40#,16#45#,16#46#,16#4f#,16#4c#,16#49#,16#4a#,
	16#6b#,16#68#,16#6d#,16#6e#,16#67#,16#64#,16#61#,16#62#,16#73#,16#70#,16#75#,16#76#,16#7f#,16#7c#,16#79#,16#7a#,
	16#3b#,16#38#,16#3d#,16#3e#,16#37#,16#34#,16#31#,16#32#,16#23#,16#20#,16#25#,16#26#,16#2f#,16#2c#,16#29#,16#2a#,
	16#0b#,16#08#,16#0d#,16#0e#,16#07#,16#04#,16#01#,16#02#,16#13#,16#10#,16#15#,16#16#,16#1f#,16#1c#,16#19#,16#1a#);

  -----------------------------------------------------------------------------
  -- Signals
  -----------------------------------------------------------------------------
  signal Matrix_D 		 : Matrix;
  signal Matrix_D_Times2 : Matrix;
  signal Matrix_D_Times3 : Matrix;
  
begin  -- architecture Behavioral
	process (Matrix_D, In_DI, Matrix_D_Times2, Matrix_D_Times3)
	begin
	for i in 0 to 3 loop
		for j in 0 to 3 loop
			Matrix_D(i)(j) <= In_DI(i)(j);
			Matrix_D_Times2(i)(j) <= std_logic_vector(to_unsigned(times2(to_integer(unsigned(In_DI(i)(j)))), 8));
			Matrix_D_Times3(i)(j) <= std_logic_vector(to_unsigned(times3(to_integer(unsigned(In_DI(i)(j)))), 8));
		end loop;
	end loop;
	end process;
	
	
  -----------------------------------------------------------------------------
  -- Output Assignment
  -----------------------------------------------------------------------------
	process (Matrix_D, In_DI, Matrix_D_Times2, Matrix_D_Times3)
	begin
	for i in 0 to 3 loop
		Out_DO(i)(0) <= Matrix_D_Times2(i)(0) xor Matrix_D_Times3(i)(1) xor Matrix_D(i)(2) xor Matrix_D(i)(3);
		Out_DO(i)(1) <= Matrix_D(i)(0) xor Matrix_D_Times2(i)(1) xor Matrix_D_Times3(i)(2) xor Matrix_D(i)(3);
		Out_DO(i)(2) <= Matrix_D(i)(0) xor Matrix_D(i)(1) xor Matrix_D_Times2(i)(2) xor Matrix_D_Times3(i)(3);
		Out_DO(i)(3) <= Matrix_D_Times3(i)(0) xor Matrix_D(i)(1) xor Matrix_D(i)(2) xor Matrix_D_Times2(i)(3);
	end loop;
	end process;
  
end architecture Behavioral;